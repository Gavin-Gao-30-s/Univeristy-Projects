library verilog;
use verilog.vl_types.all;
entity Central_RegisterFile_vlg_vec_tst is
end Central_RegisterFile_vlg_vec_tst;
