library verilog;
use verilog.vl_types.all;
entity SignleCycleProcessor_vlg_vec_tst is
end SignleCycleProcessor_vlg_vec_tst;
