library verilog;
use verilog.vl_types.all;
entity OneBitRegister_vlg_vec_tst is
end OneBitRegister_vlg_vec_tst;
