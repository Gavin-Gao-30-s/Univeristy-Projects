library verilog;
use verilog.vl_types.all;
entity ALU_12b_vlg_vec_tst is
end ALU_12b_vlg_vec_tst;
