library verilog;
use verilog.vl_types.all;
entity ALU_7bit_vlg_vec_tst is
end ALU_7bit_vlg_vec_tst;
