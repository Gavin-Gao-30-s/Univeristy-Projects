library verilog;
use verilog.vl_types.all;
entity fullAdder8_bit_plus4_vlg_sample_tst is
    port(
        A               : in     vl_logic_vector(7 downto 0);
        sampler_tx      : out    vl_logic
    );
end fullAdder8_bit_plus4_vlg_sample_tst;
