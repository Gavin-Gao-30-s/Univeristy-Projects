library verilog;
use verilog.vl_types.all;
entity fouronemux_vlg_check_tst is
    port(
        f               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end fouronemux_vlg_check_tst;
