library verilog;
use verilog.vl_types.all;
entity counter_test_vlg_vec_tst is
end counter_test_vlg_vec_tst;
