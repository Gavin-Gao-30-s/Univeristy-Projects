library verilog;
use verilog.vl_types.all;
entity fourbitcounter_vlg_vec_tst is
end fourbitcounter_vlg_vec_tst;
