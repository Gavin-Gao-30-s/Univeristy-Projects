library verilog;
use verilog.vl_types.all;
entity Extender_8to12_vlg_vec_tst is
end Extender_8to12_vlg_vec_tst;
