library verilog;
use verilog.vl_types.all;
entity bi_shift_12bit_filledWith1_vlg_vec_tst is
end bi_shift_12bit_filledWith1_vlg_vec_tst;
