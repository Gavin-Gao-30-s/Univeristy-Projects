library verilog;
use verilog.vl_types.all;
entity incrementor_7bit_vlg_vec_tst is
end incrementor_7bit_vlg_vec_tst;
