library verilog;
use verilog.vl_types.all;
entity testControlLogic_vlg_vec_tst is
end testControlLogic_vlg_vec_tst;
