library verilog;
use verilog.vl_types.all;
entity data_memory_vlg_vec_tst is
end data_memory_vlg_vec_tst;
