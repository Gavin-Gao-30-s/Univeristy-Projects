library verilog;
use verilog.vl_types.all;
entity control_logic_vlg_vec_tst is
end control_logic_vlg_vec_tst;
