library verilog;
use verilog.vl_types.all;
entity test_shiftReg2_vlg_vec_tst is
end test_shiftReg2_vlg_vec_tst;
