library verilog;
use verilog.vl_types.all;
entity test8bitConnection_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        data            : in     vl_logic_vector(7 downto 0);
        load            : in     vl_logic;
        RST             : in     vl_logic;
        shiftL          : in     vl_logic;
        shiftR          : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end test8bitConnection_vlg_sample_tst;
