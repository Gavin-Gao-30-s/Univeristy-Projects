library verilog;
use verilog.vl_types.all;
entity JumpAddress_vlg_vec_tst is
end JumpAddress_vlg_vec_tst;
