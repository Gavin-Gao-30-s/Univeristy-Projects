library verilog;
use verilog.vl_types.all;
entity data_memory_vlg_check_tst is
    port(
        read_data       : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end data_memory_vlg_check_tst;
