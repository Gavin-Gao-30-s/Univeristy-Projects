library verilog;
use verilog.vl_types.all;
entity RoundingUnit_vlg_vec_tst is
end RoundingUnit_vlg_vec_tst;
