library verilog;
use verilog.vl_types.all;
entity ID_EX_vlg_sample_tst is
    port(
        i_clock         : in     vl_logic;
        i_enable        : in     vl_logic;
        i_EX_ALUOp      : in     vl_logic_vector(1 downto 0);
        i_EX_ALUSrc     : in     vl_logic;
        i_EX_RegDst     : in     vl_logic;
        i_M_MemRead     : in     vl_logic;
        i_M_MemWrite    : in     vl_logic;
        i_Offset8       : in     vl_logic_vector(7 downto 0);
        i_Rd            : in     vl_logic_vector(2 downto 0);
        i_ReadData1     : in     vl_logic_vector(7 downto 0);
        i_ReadData2     : in     vl_logic_vector(7 downto 0);
        i_reset         : in     vl_logic;
        i_Rs            : in     vl_logic_vector(2 downto 0);
        i_Rt            : in     vl_logic_vector(2 downto 0);
        i_WB_MemToReg   : in     vl_logic;
        i_WB_RegWrite   : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end ID_EX_vlg_sample_tst;
