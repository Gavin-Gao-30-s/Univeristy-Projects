library verilog;
use verilog.vl_types.all;
entity ALU_12bit_vlg_vec_tst is
end ALU_12bit_vlg_vec_tst;
