library verilog;
use verilog.vl_types.all;
entity MUX2_5bits_vlg_vec_tst is
end MUX2_5bits_vlg_vec_tst;
