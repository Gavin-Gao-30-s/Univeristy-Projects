library verilog;
use verilog.vl_types.all;
entity incrementor_reg_vlg_vec_tst is
end incrementor_reg_vlg_vec_tst;
