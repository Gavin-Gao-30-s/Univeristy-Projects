library verilog;
use verilog.vl_types.all;
entity Down_Counter_test_vlg_vec_tst is
end Down_Counter_test_vlg_vec_tst;
