library verilog;
use verilog.vl_types.all;
entity Comparator_4bit_vlg_vec_tst is
end Comparator_4bit_vlg_vec_tst;
