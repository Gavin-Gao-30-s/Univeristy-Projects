library verilog;
use verilog.vl_types.all;
entity DifferenceChecker_vlg_vec_tst is
end DifferenceChecker_vlg_vec_tst;
