library verilog;
use verilog.vl_types.all;
entity pipeline_processor_vlg_vec_tst is
end pipeline_processor_vlg_vec_tst;
