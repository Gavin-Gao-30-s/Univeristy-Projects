library verilog;
use verilog.vl_types.all;
entity MEM_WB_vlg_vec_tst is
end MEM_WB_vlg_vec_tst;
