library verilog;
use verilog.vl_types.all;
entity Counter_4bit_vlg_vec_tst is
end Counter_4bit_vlg_vec_tst;
