library verilog;
use verilog.vl_types.all;
entity Register8bit_vlg_vec_tst is
end Register8bit_vlg_vec_tst;
