library verilog;
use verilog.vl_types.all;
entity EX_MEM_vlg_vec_tst is
end EX_MEM_vlg_vec_tst;
