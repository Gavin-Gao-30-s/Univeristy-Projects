library verilog;
use verilog.vl_types.all;
entity ID_EX_vlg_vec_tst is
end ID_EX_vlg_vec_tst;
