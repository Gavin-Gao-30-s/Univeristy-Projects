library verilog;
use verilog.vl_types.all;
entity MUX2_8bit_vlg_vec_tst is
end MUX2_8bit_vlg_vec_tst;
