library verilog;
use verilog.vl_types.all;
entity fouronemux_vlg_vec_tst is
end fouronemux_vlg_vec_tst;
