library verilog;
use verilog.vl_types.all;
entity DATAPATH is
    port(
        A_eq_B          : out    vl_logic;
        sel1            : in     vl_logic;
        expA            : in     vl_logic_vector(6 downto 0);
        expB            : in     vl_logic_vector(6 downto 0);
        Matched         : out    vl_logic;
        clk             : in     vl_logic;
        load1           : in     vl_logic;
        count1          : in     vl_logic;
        rst             : in     vl_logic;
        A_gt_B          : out    vl_logic;
        Valid           : out    vl_logic;
        Cout            : out    vl_logic;
        loadALU         : in     vl_logic;
        sel5            : in     vl_logic;
        sel3            : in     vl_logic;
        mantissaA       : in     vl_logic_vector(7 downto 0);
        mantissaB       : in     vl_logic_vector(7 downto 0);
        load2           : in     vl_logic;
        shiftR1         : in     vl_logic;
        sel4            : in     vl_logic;
        isAdd           : out    vl_logic;
        signA           : in     vl_logic;
        signB           : in     vl_logic;
        isSub           : out    vl_logic;
        normalized      : out    vl_logic;
        shiftRMAN       : out    vl_logic;
        signOut         : out    vl_logic;
        absDiffofExp    : out    vl_logic_vector(3 downto 0);
        ALU_Result      : out    vl_logic_vector(11 downto 0);
        Counter_out     : out    vl_logic_vector(3 downto 0);
        DFC_out         : out    vl_logic_vector(3 downto 0);
        expOut          : out    vl_logic_vector(6 downto 0);
        Round           : in     vl_logic;
        DEC             : in     vl_logic;
        INC             : in     vl_logic;
        load4           : in     vl_logic;
        sel2            : in     vl_logic;
        load3           : in     vl_logic;
        shiftL          : in     vl_logic;
        shiftR2         : in     vl_logic;
        Extender_out    : out    vl_logic_vector(11 downto 0);
        incrementor_out : out    vl_logic_vector(6 downto 0);
        mantissaOut     : out    vl_logic_vector(7 downto 0);
        shiftReg2_out   : out    vl_logic_vector(11 downto 0);
        shiftReg_out    : out    vl_logic_vector(11 downto 0)
    );
end DATAPATH;
