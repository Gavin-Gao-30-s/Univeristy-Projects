library verilog;
use verilog.vl_types.all;
entity Incrementor_vlg_vec_tst is
end Incrementor_vlg_vec_tst;
