library verilog;
use verilog.vl_types.all;
entity test8bitConnection_vlg_check_tst is
    port(
        \out\           : in     vl_logic_vector(11 downto 0);
        sampler_rx      : in     vl_logic
    );
end test8bitConnection_vlg_check_tst;
