LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_arith.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY instruction_memory IS
    PORT (
        address  : IN  std_logic_vector(7 DOWNTO 0); -- 8-bit address for 256 locations
        instruction : OUT std_logic_vector(31 DOWNTO 0)
    );
END instruction_memory;

ARCHITECTURE rtl OF instruction_memory IS
    TYPE rom_type IS ARRAY (0 TO 255) OF std_logic_vector(31 DOWNTO 0);
    
    CONSTANT rom : rom_type := (
     -- Address 00 (0x00): lw $2, 0($0) ; Load value from memory(00) -> $t2 = 55
        0  => X"8C020000",  
        -- Address 04 (0x04): lw $3, 1($0) ; Load value from memory(01) -> $t3 = AA
        4  => X"8C030001",  
        -- Address 08 (0x08): sub $1, $3, $2 ; $t1 = $t3 - $t2 = AA - 55 = 55 (Fixed)
        8  => X"00620822",  
        -- Address 12 (0x0C): or $4, $1, $3 ; $t4 = $t1 OR $t3 = 55 OR AA = FF
        12 => X"00232025",  
        -- Address 16 (0x10): sw $4, 3($0) ; Store $t4 (FF) into memory(03)
        16 => X"AC040003",  
        -- Address 20 (0x14): add $1, $2, $3 ; $t1 = $t2 + $t3 = 55 + AA = FF
        20 => X"00430820",  
        -- Address 24 (0x18): sw $1, 4($0) ; Store $t1 (FF) into memory(04)
        24 => X"AC010004",  
        -- Address 28 (0x1C): lw $2, 3($0) ; Load memory(03) -> $t2 = FF
        28 => X"8C020003",  
        -- Address 32 (0x20): lw $3, 4($0) ; Load memory(04) -> $t3 = FF
        32 => X"8C030004",  
        -- Address 36 (0x24): j 11 ; Jump to address 44 (0x2C)
        36 => X"0800000B",  
        -- Address 40 (0x28): beq $1, $2, -8 ; Test if $t1 == $t2 (FF == FF?)
        40 => X"1022FFFD",  
        -- Address 44 (0x2C):  beq $1, $1, -44 ; Loop back to beginning if $t1 == $t1
        44 => X"1021FFF4",  
        
        -- Fill remaining with NOP (00000000)
        OTHERS => X"00000000"
    );
BEGIN
    instruction <= rom(CONV_INTEGER(address));
END rtl;

