library verilog;
use verilog.vl_types.all;
entity Incrementor_7Bit_vlg_vec_tst is
end Incrementor_7Bit_vlg_vec_tst;
