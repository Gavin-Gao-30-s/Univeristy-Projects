library verilog;
use verilog.vl_types.all;
entity MUX4to1_vlg_vec_tst is
end MUX4to1_vlg_vec_tst;
