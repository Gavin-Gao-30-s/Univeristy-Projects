library verilog;
use verilog.vl_types.all;
entity ALU_With_Shift_vlg_vec_tst is
end ALU_With_Shift_vlg_vec_tst;
