library verilog;
use verilog.vl_types.all;
entity fullAdder8_bit_plus4_vlg_vec_tst is
end fullAdder8_bit_plus4_vlg_vec_tst;
