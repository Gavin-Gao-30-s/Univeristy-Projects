library verilog;
use verilog.vl_types.all;
entity bi_shift_12bit_vlg_check_tst is
    port(
        O_0             : in     vl_logic;
        O_1             : in     vl_logic;
        O_2             : in     vl_logic;
        O_3             : in     vl_logic;
        O_4             : in     vl_logic;
        O_5             : in     vl_logic;
        O_6             : in     vl_logic;
        O_7             : in     vl_logic;
        O_8             : in     vl_logic;
        O_9             : in     vl_logic;
        O_10            : in     vl_logic;
        O_11            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end bi_shift_12bit_vlg_check_tst;
