library verilog;
use verilog.vl_types.all;
entity FP_16bit_Adder_vlg_vec_tst is
end FP_16bit_Adder_vlg_vec_tst;
