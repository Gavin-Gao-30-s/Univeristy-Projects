library verilog;
use verilog.vl_types.all;
entity Shift_4bit_test_vlg_check_tst is
    port(
        O_0             : in     vl_logic;
        O_1             : in     vl_logic;
        O_2             : in     vl_logic;
        O_3             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Shift_4bit_test_vlg_check_tst;
