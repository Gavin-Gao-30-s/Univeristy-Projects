library verilog;
use verilog.vl_types.all;
entity test8bitConnection_vlg_vec_tst is
end test8bitConnection_vlg_vec_tst;
