library verilog;
use verilog.vl_types.all;
entity ALU_8bit_vlg_vec_tst is
end ALU_8bit_vlg_vec_tst;
