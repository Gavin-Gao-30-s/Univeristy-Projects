library verilog;
use verilog.vl_types.all;
entity Comparator_7bit_vlg_vec_tst is
end Comparator_7bit_vlg_vec_tst;
