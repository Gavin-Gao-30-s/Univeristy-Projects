library verilog;
use verilog.vl_types.all;
entity IF_ID_vlg_vec_tst is
end IF_ID_vlg_vec_tst;
