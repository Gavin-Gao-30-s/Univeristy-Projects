library verilog;
use verilog.vl_types.all;
entity debouncer_2_vlg_vec_tst is
end debouncer_2_vlg_vec_tst;
