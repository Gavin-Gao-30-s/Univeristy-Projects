library verilog;
use verilog.vl_types.all;
entity Shift_4bit_test_vlg_vec_tst is
end Shift_4bit_test_vlg_vec_tst;
