library verilog;
use verilog.vl_types.all;
entity enabledSRLatch_vlg_vec_tst is
end enabledSRLatch_vlg_vec_tst;
