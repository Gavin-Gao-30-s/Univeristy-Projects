library verilog;
use verilog.vl_types.all;
entity instruction_memory_vlg_vec_tst is
end instruction_memory_vlg_vec_tst;
